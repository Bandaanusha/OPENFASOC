MACRO VCO
  ORIGIN 0 0 ;
  FOREIGN VCO 0 0 ;
  SIZE 15.48 BY 30.24 ;
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
      LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
      LAYER M3 ;
        RECT 11.04 11.155 11.32 11.525 ;
      LAYER M2 ;
        RECT 9.46 11.2 11.18 11.48 ;
      LAYER M3 ;
        RECT 9.32 11.155 9.6 11.525 ;
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
      LAYER M3 ;
        RECT 9.32 11.155 9.6 11.525 ;
      LAYER M4 ;
        RECT 4.3 10.94 9.46 11.74 ;
      LAYER M3 ;
        RECT 4.16 11.155 4.44 11.525 ;
      LAYER M4 ;
        RECT 6.715 10.94 7.045 11.74 ;
      LAYER M3 ;
        RECT 6.74 11.155 7.02 11.525 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
      LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
      LAYER M3 ;
        RECT 11.04 3.595 11.32 3.965 ;
      LAYER M2 ;
        RECT 9.46 3.64 11.18 3.92 ;
      LAYER M3 ;
        RECT 9.32 3.595 9.6 3.965 ;
      LAYER M3 ;
        RECT 6.31 0.68 6.59 6.46 ;
      LAYER M3 ;
        RECT 9.32 3.175 9.6 3.545 ;
      LAYER M2 ;
        RECT 6.45 3.22 9.46 3.5 ;
      LAYER M3 ;
        RECT 6.31 3.175 6.59 3.545 ;
    END
  END VDD
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
      LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
      LAYER M2 ;
        RECT 8.44 7.84 8.76 8.12 ;
      LAYER M3 ;
        RECT 8.46 7.14 8.74 7.98 ;
      LAYER M2 ;
        RECT 8.44 7 8.76 7.28 ;
    END
  END OUT
  PIN IN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
      LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
      LAYER M2 ;
        RECT 3.87 12.04 5.59 12.32 ;
    END
  END IN
  OBS 
  LAYER M3 ;
        RECT 4.16 23.36 4.44 29.56 ;
  LAYER M3 ;
        RECT 5.88 23.36 6.16 29.56 ;
  LAYER M3 ;
        RECT 4.16 26.275 4.44 26.645 ;
  LAYER M2 ;
        RECT 4.3 26.32 6.02 26.6 ;
  LAYER M3 ;
        RECT 5.88 26.275 6.16 26.645 ;
  LAYER M3 ;
        RECT 13.62 23.36 13.9 29.56 ;
  LAYER M3 ;
        RECT 13.62 8.24 13.9 14.44 ;
  LAYER M3 ;
        RECT 13.62 22.68 13.9 23.52 ;
  LAYER M2 ;
        RECT 13.33 22.54 13.76 22.82 ;
  LAYER M1 ;
        RECT 13.205 15.12 13.455 22.68 ;
  LAYER M2 ;
        RECT 13.33 14.98 13.76 15.26 ;
  LAYER M3 ;
        RECT 13.62 14.28 13.9 15.12 ;
  LAYER M3 ;
        RECT 11.04 23.36 11.32 29.56 ;
  LAYER M3 ;
        RECT 9.32 23.36 9.6 29.56 ;
  LAYER M3 ;
        RECT 11.04 26.275 11.32 26.645 ;
  LAYER M2 ;
        RECT 9.46 26.32 11.18 26.6 ;
  LAYER M3 ;
        RECT 9.32 26.275 9.6 26.645 ;
  LAYER M3 ;
        RECT 0.72 19.16 1 25.36 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M3 ;
        RECT 5.88 25.855 6.16 26.225 ;
  LAYER M2 ;
        RECT 6.02 25.9 13.76 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.855 13.9 26.225 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.855 9.6 26.225 ;
  LAYER M3 ;
        RECT 4.16 23.755 4.44 24.125 ;
  LAYER M2 ;
        RECT 0.86 23.8 4.3 24.08 ;
  LAYER M3 ;
        RECT 0.72 23.755 1 24.125 ;
  LAYER M3 ;
        RECT 13.62 8.635 13.9 9.005 ;
  LAYER M2 ;
        RECT 4.73 8.68 13.76 8.96 ;
  LAYER M1 ;
        RECT 4.605 7.98 4.855 8.82 ;
  LAYER M2 ;
        RECT 3.87 7.84 4.73 8.12 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M2 ;
        RECT 0.7 23.8 1.02 24.08 ;
  LAYER M3 ;
        RECT 0.72 23.78 1 24.1 ;
  LAYER M2 ;
        RECT 4.14 23.8 4.46 24.08 ;
  LAYER M3 ;
        RECT 4.16 23.78 4.44 24.1 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M2 ;
        RECT 0.7 23.8 1.02 24.08 ;
  LAYER M3 ;
        RECT 0.72 23.78 1 24.1 ;
  LAYER M2 ;
        RECT 4.14 23.8 4.46 24.08 ;
  LAYER M3 ;
        RECT 4.16 23.78 4.44 24.1 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 8.735 4.855 8.905 ;
  LAYER M2 ;
        RECT 4.56 8.68 4.9 8.96 ;
  LAYER M2 ;
        RECT 0.7 23.8 1.02 24.08 ;
  LAYER M3 ;
        RECT 0.72 23.78 1 24.1 ;
  LAYER M2 ;
        RECT 4.14 23.8 4.46 24.08 ;
  LAYER M3 ;
        RECT 4.16 23.78 4.44 24.1 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 8.68 13.92 8.96 ;
  LAYER M3 ;
        RECT 13.62 8.66 13.9 8.98 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 8.735 4.855 8.905 ;
  LAYER M2 ;
        RECT 4.56 8.68 4.9 8.96 ;
  LAYER M2 ;
        RECT 0.7 23.8 1.02 24.08 ;
  LAYER M3 ;
        RECT 0.72 23.78 1 24.1 ;
  LAYER M2 ;
        RECT 4.14 23.8 4.46 24.08 ;
  LAYER M3 ;
        RECT 4.16 23.78 4.44 24.1 ;
  LAYER M2 ;
        RECT 5.86 25.9 6.18 26.18 ;
  LAYER M3 ;
        RECT 5.88 25.88 6.16 26.2 ;
  LAYER M2 ;
        RECT 9.3 25.9 9.62 26.18 ;
  LAYER M3 ;
        RECT 9.32 25.88 9.6 26.2 ;
  LAYER M2 ;
        RECT 13.6 8.68 13.92 8.96 ;
  LAYER M3 ;
        RECT 13.62 8.66 13.9 8.98 ;
  LAYER M2 ;
        RECT 13.6 25.9 13.92 26.18 ;
  LAYER M3 ;
        RECT 13.62 25.88 13.9 26.2 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M3 ;
        RECT 5.88 15.8 6.16 22 ;
  LAYER M3 ;
        RECT 4.16 18.715 4.44 19.085 ;
  LAYER M2 ;
        RECT 4.3 18.76 6.02 19.04 ;
  LAYER M3 ;
        RECT 5.88 18.715 6.16 19.085 ;
  LAYER M3 ;
        RECT 13.62 15.8 13.9 22 ;
  LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
  LAYER M3 ;
        RECT 13.62 16.195 13.9 16.565 ;
  LAYER M2 ;
        RECT 13.33 16.24 13.76 16.52 ;
  LAYER M3 ;
        RECT 13.19 7.56 13.47 16.38 ;
  LAYER M2 ;
        RECT 13.33 7.42 13.76 7.7 ;
  LAYER M3 ;
        RECT 13.62 6.72 13.9 7.56 ;
  LAYER M3 ;
        RECT 11.04 15.8 11.32 22 ;
  LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
  LAYER M3 ;
        RECT 11.04 18.715 11.32 19.085 ;
  LAYER M2 ;
        RECT 9.46 18.76 11.18 19.04 ;
  LAYER M3 ;
        RECT 9.32 18.715 9.6 19.085 ;
  LAYER M2 ;
        RECT 5.42 6.58 6.62 6.86 ;
  LAYER M3 ;
        RECT 0.72 11.6 1 17.8 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 6.02 15.98 13.33 16.78 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M4 ;
        RECT 7.74 7.16 13.33 7.96 ;
  LAYER M3 ;
        RECT 7.6 6.72 7.88 7.56 ;
  LAYER M2 ;
        RECT 6.45 6.58 7.74 6.86 ;
  LAYER M3 ;
        RECT 4.16 16.195 4.44 16.565 ;
  LAYER M2 ;
        RECT 0.86 16.24 4.3 16.52 ;
  LAYER M3 ;
        RECT 0.72 16.195 1 16.565 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 7.6 7.375 7.88 7.745 ;
  LAYER M4 ;
        RECT 7.575 7.16 7.905 7.96 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M4 ;
        RECT 13.165 7.16 13.495 7.96 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 7.6 7.375 7.88 7.745 ;
  LAYER M4 ;
        RECT 7.575 7.16 7.905 7.96 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M4 ;
        RECT 13.165 7.16 13.495 7.96 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M2 ;
        RECT 0.7 16.24 1.02 16.52 ;
  LAYER M3 ;
        RECT 0.72 16.22 1 16.54 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 7.6 7.375 7.88 7.745 ;
  LAYER M4 ;
        RECT 7.575 7.16 7.905 7.96 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M4 ;
        RECT 13.165 7.16 13.495 7.96 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M2 ;
        RECT 0.7 16.24 1.02 16.52 ;
  LAYER M3 ;
        RECT 0.72 16.22 1 16.54 ;
  LAYER M2 ;
        RECT 4.14 16.24 4.46 16.52 ;
  LAYER M3 ;
        RECT 4.16 16.22 4.44 16.54 ;
  LAYER M2 ;
        RECT 7.58 6.58 7.9 6.86 ;
  LAYER M3 ;
        RECT 7.6 6.56 7.88 6.88 ;
  LAYER M3 ;
        RECT 5.88 16.195 6.16 16.565 ;
  LAYER M4 ;
        RECT 5.855 15.98 6.185 16.78 ;
  LAYER M3 ;
        RECT 7.6 7.375 7.88 7.745 ;
  LAYER M4 ;
        RECT 7.575 7.16 7.905 7.96 ;
  LAYER M3 ;
        RECT 9.32 16.195 9.6 16.565 ;
  LAYER M4 ;
        RECT 9.295 15.98 9.625 16.78 ;
  LAYER M3 ;
        RECT 13.19 7.375 13.47 7.745 ;
  LAYER M4 ;
        RECT 13.165 7.16 13.495 7.96 ;
  LAYER M3 ;
        RECT 13.19 16.195 13.47 16.565 ;
  LAYER M4 ;
        RECT 13.165 15.98 13.495 16.78 ;
  LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
  LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
  LAYER M2 ;
        RECT 2.85 27.16 3.17 27.44 ;
  LAYER M1 ;
        RECT 2.885 18.06 3.135 27.3 ;
  LAYER M2 ;
        RECT 2.85 17.92 3.17 18.2 ;
  LAYER M2 ;
        RECT 1.12 18.76 2.32 19.04 ;
  LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
  LAYER M2 ;
        RECT 1.56 18.76 1.88 19.04 ;
  LAYER M3 ;
        RECT 1.58 18.06 1.86 18.9 ;
  LAYER M2 ;
        RECT 1.56 17.92 1.88 18.2 ;
  LAYER M1 ;
        RECT 2.885 18.815 3.135 18.985 ;
  LAYER M2 ;
        RECT 2.15 18.76 3.01 19.04 ;
  LAYER M1 ;
        RECT 2.885 18.815 3.135 18.985 ;
  LAYER M2 ;
        RECT 2.84 18.76 3.18 19.04 ;
  LAYER M1 ;
        RECT 2.885 18.815 3.135 18.985 ;
  LAYER M2 ;
        RECT 2.84 18.76 3.18 19.04 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M2 ;
        RECT 6.28 22.12 7.48 22.4 ;
  LAYER M2 ;
        RECT 6.72 22.96 7.04 23.24 ;
  LAYER M3 ;
        RECT 6.74 22.26 7.02 23.1 ;
  LAYER M2 ;
        RECT 6.72 22.12 7.04 22.4 ;
  LAYER M2 ;
        RECT 14.02 27.16 15.22 27.44 ;
  LAYER M2 ;
        RECT 14.02 17.92 15.22 18.2 ;
  LAYER M2 ;
        RECT 14.03 27.16 14.35 27.44 ;
  LAYER M3 ;
        RECT 14.05 18.06 14.33 27.3 ;
  LAYER M2 ;
        RECT 14.03 17.92 14.35 18.2 ;
  LAYER M3 ;
        RECT 6.74 22.495 7.02 22.865 ;
  LAYER M4 ;
        RECT 6.88 22.28 14.19 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.495 14.33 22.865 ;
  LAYER M3 ;
        RECT 6.74 22.495 7.02 22.865 ;
  LAYER M4 ;
        RECT 6.715 22.28 7.045 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.495 14.33 22.865 ;
  LAYER M4 ;
        RECT 14.025 22.28 14.355 23.08 ;
  LAYER M3 ;
        RECT 6.74 22.495 7.02 22.865 ;
  LAYER M4 ;
        RECT 6.715 22.28 7.045 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.495 14.33 22.865 ;
  LAYER M4 ;
        RECT 14.025 22.28 14.355 23.08 ;
  LAYER M2 ;
        RECT 14.02 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 14.02 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.14 14.76 7.98 ;
  LAYER M2 ;
        RECT 14.46 7 14.78 7.28 ;
  LAYER M2 ;
        RECT 11.44 27.16 12.64 27.44 ;
  LAYER M2 ;
        RECT 11.44 17.92 12.64 18.2 ;
  LAYER M2 ;
        RECT 11.45 27.16 11.77 27.44 ;
  LAYER M3 ;
        RECT 11.47 18.06 11.75 27.3 ;
  LAYER M2 ;
        RECT 11.45 17.92 11.77 18.2 ;
  LAYER M2 ;
        RECT 11.44 12.04 12.64 12.32 ;
  LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
  LAYER M2 ;
        RECT 11.45 12.04 11.77 12.32 ;
  LAYER M3 ;
        RECT 11.47 2.94 11.75 12.18 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M2 ;
        RECT 13.33 7.84 14.19 8.12 ;
  LAYER M1 ;
        RECT 13.205 7.98 13.455 9.24 ;
  LAYER M2 ;
        RECT 12.9 9.1 13.33 9.38 ;
  LAYER M1 ;
        RECT 12.775 9.24 13.025 18.06 ;
  LAYER M2 ;
        RECT 12.47 17.92 12.9 18.2 ;
  LAYER M1 ;
        RECT 12.775 12.095 13.025 12.265 ;
  LAYER M2 ;
        RECT 12.47 12.04 12.9 12.32 ;
  LAYER M1 ;
        RECT 12.775 9.155 13.025 9.325 ;
  LAYER M2 ;
        RECT 12.73 9.1 13.07 9.38 ;
  LAYER M1 ;
        RECT 12.775 17.975 13.025 18.145 ;
  LAYER M2 ;
        RECT 12.73 17.92 13.07 18.2 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.065 ;
  LAYER M2 ;
        RECT 13.16 7.84 13.5 8.12 ;
  LAYER M1 ;
        RECT 13.205 9.155 13.455 9.325 ;
  LAYER M2 ;
        RECT 13.16 9.1 13.5 9.38 ;
  LAYER M1 ;
        RECT 12.775 9.155 13.025 9.325 ;
  LAYER M2 ;
        RECT 12.73 9.1 13.07 9.38 ;
  LAYER M1 ;
        RECT 12.775 17.975 13.025 18.145 ;
  LAYER M2 ;
        RECT 12.73 17.92 13.07 18.2 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.065 ;
  LAYER M2 ;
        RECT 13.16 7.84 13.5 8.12 ;
  LAYER M1 ;
        RECT 13.205 9.155 13.455 9.325 ;
  LAYER M2 ;
        RECT 13.16 9.1 13.5 9.38 ;
  LAYER M1 ;
        RECT 12.775 9.155 13.025 9.325 ;
  LAYER M2 ;
        RECT 12.73 9.1 13.07 9.38 ;
  LAYER M1 ;
        RECT 12.775 12.095 13.025 12.265 ;
  LAYER M2 ;
        RECT 12.73 12.04 13.07 12.32 ;
  LAYER M1 ;
        RECT 12.775 17.975 13.025 18.145 ;
  LAYER M2 ;
        RECT 12.73 17.92 13.07 18.2 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.065 ;
  LAYER M2 ;
        RECT 13.16 7.84 13.5 8.12 ;
  LAYER M1 ;
        RECT 13.205 9.155 13.455 9.325 ;
  LAYER M2 ;
        RECT 13.16 9.1 13.5 9.38 ;
  LAYER M1 ;
        RECT 12.775 9.155 13.025 9.325 ;
  LAYER M2 ;
        RECT 12.73 9.1 13.07 9.38 ;
  LAYER M1 ;
        RECT 12.775 12.095 13.025 12.265 ;
  LAYER M2 ;
        RECT 12.73 12.04 13.07 12.32 ;
  LAYER M1 ;
        RECT 12.775 17.975 13.025 18.145 ;
  LAYER M2 ;
        RECT 12.73 17.92 13.07 18.2 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.065 ;
  LAYER M2 ;
        RECT 13.16 7.84 13.5 8.12 ;
  LAYER M1 ;
        RECT 13.205 9.155 13.455 9.325 ;
  LAYER M2 ;
        RECT 13.16 9.1 13.5 9.38 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M2 ;
        RECT 8 22.12 9.2 22.4 ;
  LAYER M2 ;
        RECT 8.44 22.96 8.76 23.24 ;
  LAYER M3 ;
        RECT 8.46 22.26 8.74 23.1 ;
  LAYER M2 ;
        RECT 8.44 22.12 8.76 22.4 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 1.12 13.72 2.32 14 ;
  LAYER M2 ;
        RECT 1.13 22.96 1.45 23.24 ;
  LAYER M3 ;
        RECT 1.15 13.86 1.43 23.1 ;
  LAYER M2 ;
        RECT 1.13 13.72 1.45 14 ;
  LAYER M2 ;
        RECT 8.01 22.12 8.33 22.4 ;
  LAYER M3 ;
        RECT 8.03 21.42 8.31 22.26 ;
  LAYER M2 ;
        RECT 1.29 21.28 8.17 21.56 ;
  LAYER M3 ;
        RECT 1.15 21.235 1.43 21.605 ;
  LAYER M2 ;
        RECT 1.13 21.28 1.45 21.56 ;
  LAYER M3 ;
        RECT 1.15 21.26 1.43 21.58 ;
  LAYER M2 ;
        RECT 8.01 21.28 8.33 21.56 ;
  LAYER M3 ;
        RECT 8.03 21.26 8.31 21.58 ;
  LAYER M2 ;
        RECT 8.01 22.12 8.33 22.4 ;
  LAYER M3 ;
        RECT 8.03 22.1 8.31 22.42 ;
  LAYER M2 ;
        RECT 1.13 21.28 1.45 21.56 ;
  LAYER M3 ;
        RECT 1.15 21.26 1.43 21.58 ;
  LAYER M2 ;
        RECT 8.01 21.28 8.33 21.56 ;
  LAYER M3 ;
        RECT 8.03 21.26 8.31 21.58 ;
  LAYER M2 ;
        RECT 8.01 22.12 8.33 22.4 ;
  LAYER M3 ;
        RECT 8.03 22.1 8.31 22.42 ;
  LAYER M3 ;
        RECT 5.45 2.78 5.73 7.3 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M3 ;
        RECT 5.45 7.14 5.73 7.98 ;
  LAYER M2 ;
        RECT 5.43 7.84 5.75 8.12 ;
  LAYER M2 ;
        RECT 5.43 7.84 5.75 8.12 ;
  LAYER M3 ;
        RECT 5.45 7.82 5.73 8.14 ;
  LAYER M2 ;
        RECT 5.43 7.84 5.75 8.12 ;
  LAYER M3 ;
        RECT 5.45 7.82 5.73 8.14 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 2.84 22.12 4.04 22.4 ;
  LAYER M2 ;
        RECT 3.28 22.96 3.6 23.24 ;
  LAYER M3 ;
        RECT 3.3 22.26 3.58 23.1 ;
  LAYER M2 ;
        RECT 3.28 22.12 3.6 22.4 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M2 ;
        RECT 6.28 17.92 7.48 18.2 ;
  LAYER M2 ;
        RECT 6.29 27.16 6.61 27.44 ;
  LAYER M3 ;
        RECT 6.31 18.06 6.59 27.3 ;
  LAYER M2 ;
        RECT 6.29 17.92 6.61 18.2 ;
  LAYER M3 ;
        RECT 3.3 22.495 3.58 22.865 ;
  LAYER M2 ;
        RECT 3.44 22.54 6.45 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.495 6.59 22.865 ;
  LAYER M2 ;
        RECT 3.28 22.54 3.6 22.82 ;
  LAYER M3 ;
        RECT 3.3 22.52 3.58 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M2 ;
        RECT 3.28 22.54 3.6 22.82 ;
  LAYER M3 ;
        RECT 3.3 22.52 3.58 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 26.795 3.995 27.805 ;
  LAYER M1 ;
        RECT 3.745 28.895 3.995 29.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M2 ;
        RECT 3.27 29.26 4.47 29.54 ;
  LAYER M2 ;
        RECT 3.27 23.38 4.47 23.66 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
  LAYER M3 ;
        RECT 4.16 23.36 4.44 29.56 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 16.465 ;
  LAYER M1 ;
        RECT 3.315 18.815 3.565 22.345 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M2 ;
        RECT 3.27 15.82 4.47 16.1 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M2 ;
        RECT 2.84 22.12 4.04 22.4 ;
  LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 6.325 26.795 6.575 27.805 ;
  LAYER M1 ;
        RECT 6.325 28.895 6.575 29.905 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M2 ;
        RECT 5.85 29.26 7.05 29.54 ;
  LAYER M2 ;
        RECT 5.85 23.38 7.05 23.66 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M3 ;
        RECT 5.88 23.36 6.16 29.56 ;
  LAYER M1 ;
        RECT 6.325 18.815 6.575 22.345 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 16.465 ;
  LAYER M1 ;
        RECT 6.755 18.815 7.005 22.345 ;
  LAYER M1 ;
        RECT 5.895 18.815 6.145 22.345 ;
  LAYER M2 ;
        RECT 5.85 15.82 7.05 16.1 ;
  LAYER M2 ;
        RECT 5.85 21.7 7.05 21.98 ;
  LAYER M2 ;
        RECT 6.28 22.12 7.48 22.4 ;
  LAYER M2 ;
        RECT 6.28 17.92 7.48 18.2 ;
  LAYER M3 ;
        RECT 5.88 15.8 6.16 22 ;
  LAYER M2 ;
        RECT 14.02 22.96 15.22 23.24 ;
  LAYER M2 ;
        RECT 14.02 22.12 15.22 22.4 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.26 14.76 23.1 ;
  LAYER M2 ;
        RECT 14.46 22.12 14.78 22.4 ;
  LAYER M2 ;
        RECT 14.02 12.04 15.22 12.32 ;
  LAYER M2 ;
        RECT 14.02 2.8 15.22 3.08 ;
  LAYER M2 ;
        RECT 14.03 12.04 14.35 12.32 ;
  LAYER M3 ;
        RECT 14.05 2.94 14.33 12.18 ;
  LAYER M2 ;
        RECT 14.03 2.8 14.35 3.08 ;
  LAYER M2 ;
        RECT 14.89 22.12 15.21 22.4 ;
  LAYER M1 ;
        RECT 14.925 12.18 15.175 22.26 ;
  LAYER M2 ;
        RECT 14.89 12.04 15.21 12.32 ;
  LAYER M1 ;
        RECT 14.925 12.095 15.175 12.265 ;
  LAYER M2 ;
        RECT 14.88 12.04 15.22 12.32 ;
  LAYER M1 ;
        RECT 14.925 22.175 15.175 22.345 ;
  LAYER M2 ;
        RECT 14.88 22.12 15.22 22.4 ;
  LAYER M1 ;
        RECT 14.925 12.095 15.175 12.265 ;
  LAYER M2 ;
        RECT 14.88 12.04 15.22 12.32 ;
  LAYER M1 ;
        RECT 14.925 22.175 15.175 22.345 ;
  LAYER M2 ;
        RECT 14.88 22.12 15.22 22.4 ;
  LAYER M1 ;
        RECT 14.065 23.015 14.315 26.545 ;
  LAYER M1 ;
        RECT 14.065 26.795 14.315 27.805 ;
  LAYER M1 ;
        RECT 14.065 28.895 14.315 29.905 ;
  LAYER M1 ;
        RECT 14.495 23.015 14.745 26.545 ;
  LAYER M1 ;
        RECT 13.635 23.015 13.885 26.545 ;
  LAYER M2 ;
        RECT 13.59 29.26 14.79 29.54 ;
  LAYER M2 ;
        RECT 13.59 23.38 14.79 23.66 ;
  LAYER M2 ;
        RECT 14.02 22.96 15.22 23.24 ;
  LAYER M2 ;
        RECT 14.02 27.16 15.22 27.44 ;
  LAYER M3 ;
        RECT 13.62 23.36 13.9 29.56 ;
  LAYER M1 ;
        RECT 14.065 18.815 14.315 22.345 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 15.455 14.315 16.465 ;
  LAYER M1 ;
        RECT 14.495 18.815 14.745 22.345 ;
  LAYER M1 ;
        RECT 13.635 18.815 13.885 22.345 ;
  LAYER M2 ;
        RECT 13.59 15.82 14.79 16.1 ;
  LAYER M2 ;
        RECT 13.59 21.7 14.79 21.98 ;
  LAYER M2 ;
        RECT 14.02 22.12 15.22 22.4 ;
  LAYER M2 ;
        RECT 14.02 17.92 15.22 18.2 ;
  LAYER M3 ;
        RECT 13.62 15.8 13.9 22 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M2 ;
        RECT 13.59 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 13.59 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 14.02 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 14.02 12.04 15.22 12.32 ;
  LAYER M3 ;
        RECT 13.62 8.24 13.9 14.44 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M2 ;
        RECT 13.59 0.7 14.79 0.98 ;
  LAYER M2 ;
        RECT 13.59 6.58 14.79 6.86 ;
  LAYER M2 ;
        RECT 14.02 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 14.02 2.8 15.22 3.08 ;
  LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
  LAYER M2 ;
        RECT 11.44 22.96 12.64 23.24 ;
  LAYER M2 ;
        RECT 11.44 22.12 12.64 22.4 ;
  LAYER M2 ;
        RECT 11.88 22.96 12.2 23.24 ;
  LAYER M3 ;
        RECT 11.9 22.26 12.18 23.1 ;
  LAYER M2 ;
        RECT 11.88 22.12 12.2 22.4 ;
  LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
  LAYER M2 ;
        RECT 8 17.92 9.2 18.2 ;
  LAYER M2 ;
        RECT 8.01 27.16 8.33 27.44 ;
  LAYER M1 ;
        RECT 8.045 18.06 8.295 27.3 ;
  LAYER M2 ;
        RECT 8.01 17.92 8.33 18.2 ;
  LAYER M3 ;
        RECT 11.9 22.495 12.18 22.865 ;
  LAYER M2 ;
        RECT 8.17 22.54 12.04 22.82 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M2 ;
        RECT 8 22.54 8.34 22.82 ;
  LAYER M2 ;
        RECT 11.88 22.54 12.2 22.82 ;
  LAYER M3 ;
        RECT 11.9 22.52 12.18 22.84 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M2 ;
        RECT 8 22.54 8.34 22.82 ;
  LAYER M2 ;
        RECT 11.88 22.54 12.2 22.82 ;
  LAYER M3 ;
        RECT 11.9 22.52 12.18 22.84 ;
  LAYER M1 ;
        RECT 11.485 23.015 11.735 26.545 ;
  LAYER M1 ;
        RECT 11.485 26.795 11.735 27.805 ;
  LAYER M1 ;
        RECT 11.485 28.895 11.735 29.905 ;
  LAYER M1 ;
        RECT 11.915 23.015 12.165 26.545 ;
  LAYER M1 ;
        RECT 11.055 23.015 11.305 26.545 ;
  LAYER M2 ;
        RECT 11.01 29.26 12.21 29.54 ;
  LAYER M2 ;
        RECT 11.01 23.38 12.21 23.66 ;
  LAYER M2 ;
        RECT 11.44 22.96 12.64 23.24 ;
  LAYER M2 ;
        RECT 11.44 27.16 12.64 27.44 ;
  LAYER M3 ;
        RECT 11.04 23.36 11.32 29.56 ;
  LAYER M1 ;
        RECT 11.485 18.815 11.735 22.345 ;
  LAYER M1 ;
        RECT 11.485 17.555 11.735 18.565 ;
  LAYER M1 ;
        RECT 11.485 15.455 11.735 16.465 ;
  LAYER M1 ;
        RECT 11.915 18.815 12.165 22.345 ;
  LAYER M1 ;
        RECT 11.055 18.815 11.305 22.345 ;
  LAYER M2 ;
        RECT 11.01 15.82 12.21 16.1 ;
  LAYER M2 ;
        RECT 11.01 21.7 12.21 21.98 ;
  LAYER M2 ;
        RECT 11.44 22.12 12.64 22.4 ;
  LAYER M2 ;
        RECT 11.44 17.92 12.64 18.2 ;
  LAYER M3 ;
        RECT 11.04 15.8 11.32 22 ;
  LAYER M1 ;
        RECT 8.905 23.015 9.155 26.545 ;
  LAYER M1 ;
        RECT 8.905 26.795 9.155 27.805 ;
  LAYER M1 ;
        RECT 8.905 28.895 9.155 29.905 ;
  LAYER M1 ;
        RECT 8.475 23.015 8.725 26.545 ;
  LAYER M1 ;
        RECT 9.335 23.015 9.585 26.545 ;
  LAYER M2 ;
        RECT 8.43 29.26 9.63 29.54 ;
  LAYER M2 ;
        RECT 8.43 23.38 9.63 23.66 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
  LAYER M3 ;
        RECT 9.32 23.36 9.6 29.56 ;
  LAYER M1 ;
        RECT 8.905 18.815 9.155 22.345 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 15.455 9.155 16.465 ;
  LAYER M1 ;
        RECT 8.475 18.815 8.725 22.345 ;
  LAYER M1 ;
        RECT 9.335 18.815 9.585 22.345 ;
  LAYER M2 ;
        RECT 8.43 15.82 9.63 16.1 ;
  LAYER M2 ;
        RECT 8.43 21.7 9.63 21.98 ;
  LAYER M2 ;
        RECT 8 22.12 9.2 22.4 ;
  LAYER M2 ;
        RECT 8 17.92 9.2 18.2 ;
  LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
  LAYER M2 ;
        RECT 11.44 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 11.88 7.84 12.2 8.12 ;
  LAYER M3 ;
        RECT 11.9 7.14 12.18 7.98 ;
  LAYER M2 ;
        RECT 11.88 7 12.2 7.28 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M1 ;
        RECT 8.045 2.94 8.295 12.18 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M3 ;
        RECT 11.9 7.375 12.18 7.745 ;
  LAYER M2 ;
        RECT 8.17 7.42 12.04 7.7 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 11.88 7.42 12.2 7.7 ;
  LAYER M3 ;
        RECT 11.9 7.4 12.18 7.72 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 11.44 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 11.44 12.04 12.64 12.32 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 11.01 0.7 12.21 0.98 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
  LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 5.42 0.7 6.62 0.98 ;
  LAYER M2 ;
        RECT 4.99 6.16 7.05 6.44 ;
  LAYER M3 ;
        RECT 5.45 2.78 5.73 7.3 ;
  LAYER M2 ;
        RECT 5.42 6.58 6.62 6.86 ;
  LAYER M3 ;
        RECT 6.31 0.68 6.59 6.46 ;
  LAYER M1 ;
        RECT 1.165 18.815 1.415 22.345 ;
  LAYER M1 ;
        RECT 1.165 22.595 1.415 23.605 ;
  LAYER M1 ;
        RECT 1.165 24.695 1.415 25.705 ;
  LAYER M1 ;
        RECT 1.595 18.815 1.845 22.345 ;
  LAYER M1 ;
        RECT 0.735 18.815 0.985 22.345 ;
  LAYER M2 ;
        RECT 0.69 25.06 1.89 25.34 ;
  LAYER M2 ;
        RECT 0.69 19.18 1.89 19.46 ;
  LAYER M2 ;
        RECT 1.12 18.76 2.32 19.04 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M3 ;
        RECT 0.72 19.16 1 25.36 ;
  LAYER M1 ;
        RECT 1.165 14.615 1.415 18.145 ;
  LAYER M1 ;
        RECT 1.165 13.355 1.415 14.365 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 12.265 ;
  LAYER M1 ;
        RECT 1.595 14.615 1.845 18.145 ;
  LAYER M1 ;
        RECT 0.735 14.615 0.985 18.145 ;
  LAYER M2 ;
        RECT 0.69 11.62 1.89 11.9 ;
  LAYER M2 ;
        RECT 0.69 17.5 1.89 17.78 ;
  LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
  LAYER M2 ;
        RECT 1.12 13.72 2.32 14 ;
  LAYER M3 ;
        RECT 0.72 11.6 1 17.8 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  END 
END VCO
